
module unsaved (
	clk_clk,
	portd_external_connection_export);	

	input		clk_clk;
	output	[7:0]	portd_external_connection_export;
endmodule
