
module unsaved (
	clk_clk,
	latx_external_connection_export,
	portx_external_connection_export);	

	input		clk_clk;
	output	[7:0]	latx_external_connection_export;
	input	[1:0]	portx_external_connection_export;
endmodule
