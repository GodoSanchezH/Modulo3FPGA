-- unsaved.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unsaved is
	port (
		clk_clk                         : in  std_logic                    := '0';             --                      clk.clk
		leds_external_connection_export : out std_logic_vector(9 downto 0);                    -- leds_external_connection.export
		sw_external_connection_export   : in  std_logic_vector(1 downto 0) := (others => '0')  --   sw_external_connection.export
	);
end entity unsaved;

architecture rtl of unsaved is
	component unsaved_LEDS is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component unsaved_LEDS;

	component unsaved_SW is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component unsaved_SW;

	component unsaved_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component unsaved_jtag_uart;

	component unsaved_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component unsaved_memory;

	component unsaved_nios2 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(17 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(17 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component unsaved_nios2;

	component unsaved_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component unsaved_sysid_qsys_0;

	component unsaved_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			nios2_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_data_master_address                 : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			nios2_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_data_master_read                    : in  std_logic                     := 'X';             -- read
			nios2_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_data_master_write                   : in  std_logic                     := 'X';             -- write
			nios2_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			nios2_instruction_master_address          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			nios2_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			nios2_instruction_master_read             : in  std_logic                     := 'X';             -- read
			nios2_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_uart_avalon_jtag_slave_address       : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write         : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read          : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect    : out std_logic;                                        -- chipselect
			LEDS_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			LEDS_s1_write                             : out std_logic;                                        -- write
			LEDS_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDS_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			LEDS_s1_chipselect                        : out std_logic;                                        -- chipselect
			memory_s1_address                         : out std_logic_vector(13 downto 0);                    -- address
			memory_s1_write                           : out std_logic;                                        -- write
			memory_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			memory_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			memory_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			memory_s1_chipselect                      : out std_logic;                                        -- chipselect
			memory_s1_clken                           : out std_logic;                                        -- clken
			nios2_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			nios2_jtag_debug_module_write             : out std_logic;                                        -- write
			nios2_jtag_debug_module_read              : out std_logic;                                        -- read
			nios2_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			nios2_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			SW_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			SW_s1_write                               : out std_logic;                                        -- write
			SW_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SW_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			SW_s1_chipselect                          : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address        : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component unsaved_mm_interconnect_0;

	component unsaved_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component unsaved_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal nios2_jtag_debug_module_reset_reset                           : std_logic;                     -- nios2:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	signal nios2_data_master_readdata                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	signal nios2_data_master_waitrequest                                 : std_logic;                     -- mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	signal nios2_data_master_debugaccess                                 : std_logic;                     -- nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	signal nios2_data_master_address                                     : std_logic_vector(17 downto 0); -- nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	signal nios2_data_master_byteenable                                  : std_logic_vector(3 downto 0);  -- nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	signal nios2_data_master_read                                        : std_logic;                     -- nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	signal nios2_data_master_write                                       : std_logic;                     -- nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	signal nios2_data_master_writedata                                   : std_logic_vector(31 downto 0); -- nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	signal nios2_instruction_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	signal nios2_instruction_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	signal nios2_instruction_master_address                              : std_logic_vector(17 downto 0); -- nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	signal nios2_instruction_master_read                                 : std_logic;                     -- nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata         : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_jtag_debug_module_readdata            : std_logic_vector(31 downto 0); -- nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_jtag_debug_module_waitrequest         : std_logic;                     -- nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_jtag_debug_module_debugaccess         : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_jtag_debug_module_address             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	signal mm_interconnect_0_nios2_jtag_debug_module_read                : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	signal mm_interconnect_0_nios2_jtag_debug_module_byteenable          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	signal mm_interconnect_0_nios2_jtag_debug_module_write               : std_logic;                     -- mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	signal mm_interconnect_0_nios2_jtag_debug_module_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	signal mm_interconnect_0_memory_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	signal mm_interconnect_0_memory_s1_readdata                          : std_logic_vector(31 downto 0); -- memory:readdata -> mm_interconnect_0:memory_s1_readdata
	signal mm_interconnect_0_memory_s1_address                           : std_logic_vector(13 downto 0); -- mm_interconnect_0:memory_s1_address -> memory:address
	signal mm_interconnect_0_memory_s1_byteenable                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	signal mm_interconnect_0_memory_s1_write                             : std_logic;                     -- mm_interconnect_0:memory_s1_write -> memory:write
	signal mm_interconnect_0_memory_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:memory_s1_writedata -> memory:writedata
	signal mm_interconnect_0_memory_s1_clken                             : std_logic;                     -- mm_interconnect_0:memory_s1_clken -> memory:clken
	signal mm_interconnect_0_leds_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	signal mm_interconnect_0_leds_s1_readdata                            : std_logic_vector(31 downto 0); -- LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	signal mm_interconnect_0_leds_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDS_s1_address -> LEDS:address
	signal mm_interconnect_0_leds_s1_write                               : std_logic;                     -- mm_interconnect_0:LEDS_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	signal mm_interconnect_0_sw_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:SW_s1_chipselect -> SW:chipselect
	signal mm_interconnect_0_sw_s1_readdata                              : std_logic_vector(31 downto 0); -- SW:readdata -> mm_interconnect_0:SW_s1_readdata
	signal mm_interconnect_0_sw_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SW_s1_address -> SW:address
	signal mm_interconnect_0_sw_s1_write                                 : std_logic;                     -- mm_interconnect_0:SW_s1_write -> mm_interconnect_0_sw_s1_write:in
	signal mm_interconnect_0_sw_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:SW_s1_writedata -> SW:writedata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- SW:irq -> irq_mapper:receiver1_irq
	signal nios2_d_irq_irq                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2:d_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, memory:reset, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [memory:reset_req, nios2:reset_req, rst_translator:reset_req_in]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_leds_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> LEDS:write_n
	signal mm_interconnect_0_sw_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_sw_s1_write:inv -> SW:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [LEDS:reset_n, SW:reset_n, jtag_uart:rst_n, nios2:reset_n, sysid_qsys_0:reset_n]

begin

	leds : component unsaved_LEDS
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_external_connection_export            -- external_connection.export
		);

	sw : component unsaved_SW
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_sw_s1_address,          --                  s1.address
			write_n    => mm_interconnect_0_sw_s1_write_ports_inv,  --                    .write_n
			writedata  => mm_interconnect_0_sw_s1_writedata,        --                    .writedata
			chipselect => mm_interconnect_0_sw_s1_chipselect,       --                    .chipselect
			readdata   => mm_interconnect_0_sw_s1_readdata,         --                    .readdata
			in_port    => sw_external_connection_export,            -- external_connection.export
			irq        => irq_mapper_receiver1_irq                  --                 irq.irq
		);

	jtag_uart : component unsaved_jtag_uart
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	memory : component unsaved_memory
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,     --       .reset_req
			freeze     => '0'                                     -- (terminated)
		);

	nios2 : component unsaved_nios2
		port map (
			clk                                   => clk_clk,                                               --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,              --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                    --                          .reset_req
			d_address                             => nios2_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_data_master_read,                                --                          .read
			d_readdata                            => nios2_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_data_master_write,                               --                          .write
			d_writedata                           => nios2_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => nios2_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                   -- custom_instruction_master.readra
		);

	sysid_qsys_0 : component unsaved_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component unsaved_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                                   --                           clk_0_clk.clk
			nios2_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- nios2_reset_n_reset_bridge_in_reset.reset
			nios2_data_master_address                 => nios2_data_master_address,                                 --                   nios2_data_master.address
			nios2_data_master_waitrequest             => nios2_data_master_waitrequest,                             --                                    .waitrequest
			nios2_data_master_byteenable              => nios2_data_master_byteenable,                              --                                    .byteenable
			nios2_data_master_read                    => nios2_data_master_read,                                    --                                    .read
			nios2_data_master_readdata                => nios2_data_master_readdata,                                --                                    .readdata
			nios2_data_master_write                   => nios2_data_master_write,                                   --                                    .write
			nios2_data_master_writedata               => nios2_data_master_writedata,                               --                                    .writedata
			nios2_data_master_debugaccess             => nios2_data_master_debugaccess,                             --                                    .debugaccess
			nios2_instruction_master_address          => nios2_instruction_master_address,                          --            nios2_instruction_master.address
			nios2_instruction_master_waitrequest      => nios2_instruction_master_waitrequest,                      --                                    .waitrequest
			nios2_instruction_master_read             => nios2_instruction_master_read,                             --                                    .read
			nios2_instruction_master_readdata         => nios2_instruction_master_readdata,                         --                                    .readdata
			jtag_uart_avalon_jtag_slave_address       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --         jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                    .write
			jtag_uart_avalon_jtag_slave_read          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                    .read
			jtag_uart_avalon_jtag_slave_readdata      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                    .readdata
			jtag_uart_avalon_jtag_slave_writedata     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                    .writedata
			jtag_uart_avalon_jtag_slave_waitrequest   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                    .chipselect
			LEDS_s1_address                           => mm_interconnect_0_leds_s1_address,                         --                             LEDS_s1.address
			LEDS_s1_write                             => mm_interconnect_0_leds_s1_write,                           --                                    .write
			LEDS_s1_readdata                          => mm_interconnect_0_leds_s1_readdata,                        --                                    .readdata
			LEDS_s1_writedata                         => mm_interconnect_0_leds_s1_writedata,                       --                                    .writedata
			LEDS_s1_chipselect                        => mm_interconnect_0_leds_s1_chipselect,                      --                                    .chipselect
			memory_s1_address                         => mm_interconnect_0_memory_s1_address,                       --                           memory_s1.address
			memory_s1_write                           => mm_interconnect_0_memory_s1_write,                         --                                    .write
			memory_s1_readdata                        => mm_interconnect_0_memory_s1_readdata,                      --                                    .readdata
			memory_s1_writedata                       => mm_interconnect_0_memory_s1_writedata,                     --                                    .writedata
			memory_s1_byteenable                      => mm_interconnect_0_memory_s1_byteenable,                    --                                    .byteenable
			memory_s1_chipselect                      => mm_interconnect_0_memory_s1_chipselect,                    --                                    .chipselect
			memory_s1_clken                           => mm_interconnect_0_memory_s1_clken,                         --                                    .clken
			nios2_jtag_debug_module_address           => mm_interconnect_0_nios2_jtag_debug_module_address,         --             nios2_jtag_debug_module.address
			nios2_jtag_debug_module_write             => mm_interconnect_0_nios2_jtag_debug_module_write,           --                                    .write
			nios2_jtag_debug_module_read              => mm_interconnect_0_nios2_jtag_debug_module_read,            --                                    .read
			nios2_jtag_debug_module_readdata          => mm_interconnect_0_nios2_jtag_debug_module_readdata,        --                                    .readdata
			nios2_jtag_debug_module_writedata         => mm_interconnect_0_nios2_jtag_debug_module_writedata,       --                                    .writedata
			nios2_jtag_debug_module_byteenable        => mm_interconnect_0_nios2_jtag_debug_module_byteenable,      --                                    .byteenable
			nios2_jtag_debug_module_waitrequest       => mm_interconnect_0_nios2_jtag_debug_module_waitrequest,     --                                    .waitrequest
			nios2_jtag_debug_module_debugaccess       => mm_interconnect_0_nios2_jtag_debug_module_debugaccess,     --                                    .debugaccess
			SW_s1_address                             => mm_interconnect_0_sw_s1_address,                           --                               SW_s1.address
			SW_s1_write                               => mm_interconnect_0_sw_s1_write,                             --                                    .write
			SW_s1_readdata                            => mm_interconnect_0_sw_s1_readdata,                          --                                    .readdata
			SW_s1_writedata                           => mm_interconnect_0_sw_s1_writedata,                         --                                    .writedata
			SW_s1_chipselect                          => mm_interconnect_0_sw_s1_chipselect,                        --                                    .chipselect
			sysid_qsys_0_control_slave_address        => mm_interconnect_0_sysid_qsys_0_control_slave_address,      --          sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata       => mm_interconnect_0_sysid_qsys_0_control_slave_readdata      --                                    .readdata
		);

	irq_mapper : component unsaved_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_d_irq_irq                 --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_jtag_debug_module_reset_reset, -- reset_in0.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,  --          .reset_req
			reset_req_in0  => '0',                                 -- (terminated)
			reset_in1      => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_sw_s1_write_ports_inv <= not mm_interconnect_0_sw_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of unsaved
