mult_inst : mult PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
